library verilog;
use verilog.vl_types.all;
entity date is
    generic(
        state0          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        state1          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        state2          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        state3          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        state4          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        state5          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        scan            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        nul             : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        data0           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        data1           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1);
        data2           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0);
        data3           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1);
        data4           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        data5           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        data6           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0);
        data7           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1);
        data8           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        data9           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1);
        data10          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        data11          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1);
        data12          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0);
        data13          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        data14          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        data15          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1);
        data16          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0);
        data17          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1);
        data18          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        data19          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1);
        data20          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0);
        data21          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1);
        data22          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        data23          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1);
        data24          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0);
        data25          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1);
        data26          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0);
        data27          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1);
        data28          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0);
        data29          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1);
        data30          : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        data31          : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1)
    );
    port(
        rst             : in     vl_logic;
        clk             : in     vl_logic;
        rw              : out    vl_logic;
        rs              : out    vl_logic;
        en              : out    vl_logic;
        data            : out    vl_logic_vector(7 downto 0);
        key1            : in     vl_logic;
        key2            : in     vl_logic;
        key3            : in     vl_logic;
        led             : out    vl_logic_vector(3 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of state0 : constant is 1;
    attribute mti_svvh_generic_type of state1 : constant is 1;
    attribute mti_svvh_generic_type of state2 : constant is 1;
    attribute mti_svvh_generic_type of state3 : constant is 1;
    attribute mti_svvh_generic_type of state4 : constant is 1;
    attribute mti_svvh_generic_type of state5 : constant is 1;
    attribute mti_svvh_generic_type of scan : constant is 1;
    attribute mti_svvh_generic_type of nul : constant is 1;
    attribute mti_svvh_generic_type of data0 : constant is 1;
    attribute mti_svvh_generic_type of data1 : constant is 1;
    attribute mti_svvh_generic_type of data2 : constant is 1;
    attribute mti_svvh_generic_type of data3 : constant is 1;
    attribute mti_svvh_generic_type of data4 : constant is 1;
    attribute mti_svvh_generic_type of data5 : constant is 1;
    attribute mti_svvh_generic_type of data6 : constant is 1;
    attribute mti_svvh_generic_type of data7 : constant is 1;
    attribute mti_svvh_generic_type of data8 : constant is 1;
    attribute mti_svvh_generic_type of data9 : constant is 1;
    attribute mti_svvh_generic_type of data10 : constant is 1;
    attribute mti_svvh_generic_type of data11 : constant is 1;
    attribute mti_svvh_generic_type of data12 : constant is 1;
    attribute mti_svvh_generic_type of data13 : constant is 1;
    attribute mti_svvh_generic_type of data14 : constant is 1;
    attribute mti_svvh_generic_type of data15 : constant is 1;
    attribute mti_svvh_generic_type of data16 : constant is 1;
    attribute mti_svvh_generic_type of data17 : constant is 1;
    attribute mti_svvh_generic_type of data18 : constant is 1;
    attribute mti_svvh_generic_type of data19 : constant is 1;
    attribute mti_svvh_generic_type of data20 : constant is 1;
    attribute mti_svvh_generic_type of data21 : constant is 1;
    attribute mti_svvh_generic_type of data22 : constant is 1;
    attribute mti_svvh_generic_type of data23 : constant is 1;
    attribute mti_svvh_generic_type of data24 : constant is 1;
    attribute mti_svvh_generic_type of data25 : constant is 1;
    attribute mti_svvh_generic_type of data26 : constant is 1;
    attribute mti_svvh_generic_type of data27 : constant is 1;
    attribute mti_svvh_generic_type of data28 : constant is 1;
    attribute mti_svvh_generic_type of data29 : constant is 1;
    attribute mti_svvh_generic_type of data30 : constant is 1;
    attribute mti_svvh_generic_type of data31 : constant is 1;
end date;
